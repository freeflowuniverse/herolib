module webdav

import freeflowuniverse.herolib.ui.console
import log

// fn add_dav_headers(mut ctx Context) bool {
// 	ctx.set_custom_header('dav', '1,2') or { return ctx.server_error(err.msg()) }
// 	ctx.set_header(.allow, 'OPTIONS, PROPFIND, MKCOL, GET, HEAD, POST, PUT, DELETE, COPY, MOVE')
// 	ctx.set_custom_header('MS-Author-Via', 'DAV') or { return ctx.server_error(err.msg()) }
// 	return true
// }
