module reprompt

import freeflowuniverse.herolib.data.paramsparser
import freeflowuniverse.herolib.data.encoderhero
import freeflowuniverse.herolib.core.pathlib
import os

// your checking & initialization code if needed
fn (mut ws RepromptWorkspace) reprompt() !string {
	//TODO: fill in template based on selection
	return ""
}
