module rhai