module mycelium
