module giteaclient

import freeflowuniverse.herolib.core.base
import freeflowuniverse.herolib.core.playbook { PlayBook }
import freeflowuniverse.herolib.ui.console

__global (
	giteaclient_global  map[string]&GiteaClient
	giteaclient_default string
)

/////////FACTORY

@[params]
pub struct ArgsGet {
pub mut:
	name string
}

fn args_get(args_ ArgsGet) ArgsGet {
	mut args := args_
	if args.name == '' {
		args.name = 'default'
	}
	return args
}

pub fn get(args_ ArgsGet) !&GiteaClient {
	mut context := base.context()!
	mut args := args_get(args_)
	mut obj := GiteaClient{
		name: args.name
	}
	if args.name !in giteaclient_global {
		if !exists(args)! {
			set(obj)!
		} else {
			heroscript := context.hero_config_get('giteaclient', args.name)!
			mut obj_ := heroscript_loads(heroscript)!
			set_in_mem(obj_)!
		}
	}
	return giteaclient_global[args.name] or {
		println(giteaclient_global)
		// bug if we get here because should be in globals
		panic('could not get config for giteaclient with name, is bug:${args.name}')
	}
}

// register the config for the future
pub fn set(o GiteaClient) ! {
	set_in_mem(o)!
	mut context := base.context()!
	heroscript := heroscript_dumps(o)!
	context.hero_config_set('giteaclient', o.name, heroscript)!
}

// does the config exists?
pub fn exists(args_ ArgsGet) !bool {
	mut context := base.context()!
	mut args := args_get(args_)
	return context.hero_config_exists('giteaclient', args.name)
}

pub fn delete(args_ ArgsGet) ! {
	mut args := args_get(args_)
	mut context := base.context()!
	context.hero_config_delete('giteaclient', args.name)!
	if args.name in giteaclient_global {
		// del giteaclient_global[args.name]
	}
}

@[params]
pub struct ArgsList {
pub mut:
	fromdb bool //will load from filesystem
}


pub fn list(args ArgsList) ![]&GiteaClient {
	
	mut res := []&GiteaClient{}
	if args.name in giteaclient_global {
		res << giteaclient_global[o.name]
	}
	return res
}

// only sets in mem, does not set as config
fn set_in_mem(o GiteaClient) ! {
	mut o2 := obj_init(o)!
	giteaclient_global[o.name] = &o2
	giteaclient_default = o.name
}

pub fn play(mut plbook PlayBook) ! {
	mut install_actions := plbook.find(filter: 'giteaclient.configure')!
	if install_actions.len > 0 {
		for install_action in install_actions {
			heroscript := install_action.heroscript()
			mut obj2 := heroscript_loads(heroscript)!
			set(obj2)!
		}
	}
}

// switch instance to be used for giteaclient
pub fn switch(name string) {
	giteaclient_default = name
}

// helpers

@[params]
pub struct DefaultConfigArgs {
	instance string = 'default'
}
