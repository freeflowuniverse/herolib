module handlers

import os
import freeflowuniverse.herolib.mcp.v_do.logger
