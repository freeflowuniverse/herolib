module installers

// import freeflowuniverse.herolib.core.pathlib
// import freeflowuniverse.herolib.develop.gittools

@[params]
pub struct UploadArgs {
pub mut:
	cmdname string
	source  string
	reset   bool
}

pub fn upload_(args_ UploadArgs) ! {
	//_ := args_
	panic('to implement')
}
