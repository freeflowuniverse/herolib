module ui

// Placeholder for heroscript-specific utilities
