module location

// https://www.geonames.org/export/codes.html
