module mcp

pub type Any = []Any
	| bool
	| int
	| map[string]Any
	| string