module processmanager

import freeflowuniverse.herolib.osal

pub struct ProcessManager {
	// pub mut:
}

pub fn new() !ProcessManager {
	mut pm := ProcessManager{}
}
