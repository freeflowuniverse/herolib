module docusaurus

import os
import freeflowuniverse.herolib.core.pathlib
import freeflowuniverse.herolib.core.texttools
import freeflowuniverse.herolib.develop.gittools
import freeflowuniverse.herolib.web.siteconfig
import freeflowuniverse.herolib.ui.console
import freeflowuniverse.herolib.osal

@[params]
pub struct DSiteGetArgs {
pub mut:
	name          string
	nameshort     string
	path          string
	url           string
	path_publish  string //default empty
	// path_build    string //default empty
	production    bool
	watch_changes bool = true
	update        bool
	open          bool
	init          bool // means create new one if needed
	deploykey     string
	// config        ?Configuration
}

pub fn (mut f DocusaurusFactory) get(args_ DSiteGetArgs) !&DocSite {
	console.print_header(' Docusaurus: ${args_.name}')
	mut args := args_

	// coderoot:"${os.home_dir()}/hero/var/publishcode"
	mut gs := gittools.new(ssh_key_path: args.deploykey)!

	if args.url.len > 0 {
		args.path = gs.get_path(url: args.url)!
	}

	if args.path.trim_space() == '' {
		args.path = os.getwd()
	}
	args.path = args.path.replace('~', os.home_dir())

	configpath:='${args.path}/cfg'
	if ! os.exists(configpath) {
		return error("can't find config file in ${configpath}")
	}

	osal.rm("${args.path}/cfg/main.json")!
	osal.rm("${args.path}/cfg/footer.json")!
	osal.rm("${args.path}/cfg/navbar.json")!
	osal.rm("${args.path}/build.sh")!
	osal.rm("${args.path}/develop.sh")!
	osal.rm("${args.path}/sync.sh")!
	osal.rm("${args.path}/.DS_Store")!

	if !os.exists('${args.path}/docs') {
		if args.init {
			// Create docs directory if it doesn't exist in template or site
			os.mkdir_all('${args.path}/docs')!
			panic("implement")
		} else {
			return error("Can't find docs dir in chosen docusaurus location: ${args.path}")
		}
	}


	mut myconfig:=config_load(configpath)!

	if myconfig.main.name.len == 0 {
		myconfig.main.name = myconfig.main.base_url.trim_space().trim('/').trim_space()
	}

	if args.name == '' {
		args.name = myconfig.main.name
	}

	if args.nameshort.len == 0 {
		args.nameshort = args.name
	}
	args.nameshort = texttools.name_fix(args.nameshort)

	if args.path_publish == ""{
		args.path_publish = "${f.path_publish}/${args.name}"
	}

	mut mysiteconfig:=*siteconfig.new(configpath)!

	mut ds := DocSite{
		name:       args.name
		url:        args.url
		path_src:   pathlib.get_dir(path: args.path, create: false)!
		path_publish: pathlib.get_dir(path:args.path_publish)!
		args:    args
		config:  myconfig
		siteconfig: mysiteconfig //comes from the heroconfig
		factory: &f
	}
	ds.check()!

	f.sites << &ds

	return &ds
}
