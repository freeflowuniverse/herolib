module blockchain

// import freeflowuniverse.herolib.core.playbook

pub struct Controller {
}

pub fn new() !Controller {
	mut c := Controller{}
	return c
}
