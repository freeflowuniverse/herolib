module ui

// Placeholder for chat-specific utilities
