module heroscript

// Placeholder for heroscript-specific utilities

