module handlers

import os
import freeflowuniverse.herolib.mcp.v_do.logger



cmd := 'v -gc none -stats -enable-globals -show-c-output -keepc -n -w -cg -o /tmp/tester.c -g -cc tcc ${fullpath}'