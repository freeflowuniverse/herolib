module chat

// Placeholder for chat-specific utilities

