module ui

// Placeholder for heroprompt-specific utilities (if needed later)
