module heroprompt
