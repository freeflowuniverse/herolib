module playcmds

import freeflowuniverse.herolib.develop.gittools
import freeflowuniverse.herolib.core.playbook { PlayBook }
import freeflowuniverse.herolib.core.base
import freeflowuniverse.herolib.ui.console

// !!context.configure
//     name:'test'
//     coderoot:...
//     interactive:true


fn play_core(mut plbook PlayBook) ! {

	// for mut action in plbook.find(filter: 'context.configure')! {
	// 	mut p := action.params
	// 	mut session := plbook.session

	// 	if p.exists('interactive') {
	// 		session.interactive = p.get_default_false('interactive')
	// 	}

	// 	if p.exists('coderoot') {
	// 		panic('implement')
	// 		// mut coderoot := p.get_path_create('coderoot')!
	// 		// mut gs := gittools.get()!
	// 	}
	// 	action.done = true
	// }

	for action_ in plbook.find(filter: 'play.*')! {
		if action_.name == 'include' {
			console.print_debug('play run:${action_}')
			mut action := *action_
			mut playrunpath := action.params.get_default('path', '')!
			if playrunpath.len == 0 {
				action.name = 'pull'
				playrunpath = gittools.get_repo_path(
						path:action.params.get_default('path', '')!
						git_url:action.params.get_default('git_url', '')!
						git_reset:action.params.get_default_false('git_reset')
						git_pull:action.params.get_default_false('git_pull')
						)!
			}
			if playrunpath.len == 0 {
				return error("can't run a heroscript didn't find url or path.")
			}
			console.print_debug('play run path:${playrunpath}')
			plbook.add(path: playrunpath)!
		}
		if action_.name == 'echo' {
			content := action_.params.get_default('content', "didn't find content")!
			console.print_header(content)
		}
	}	

	for mut action in plbook.find(filter: 'session.')! {
		mut p := action.params
		mut session := plbook.session

		//!!session.env_set key:'JWT_SHARED_KEY' val:'...'
		if p.exists('env_set') {
			mut key := p.get('key')!
			mut val := p.get('val')!
			session.env_set(key, val)!
		}

		if p.exists('env_set_once') {
			mut key := p.get('key')!
			mut val := p.get('val')!
			session.env_set_once(key, val)!
		}		

		action.done = true
	}


	// CHANGE {...} args in plbook

	println('plbook:${plbook}')

	mut context := base.context()!
	mut session := context.session_latest()!

	sitename:=session.env_get('SITENAME') or {""}

	println('session:${session}')
	println('sitename:${sitename}')

	if true{panic("dfghjkjhgfghjk")}

	// for mut action in plbook.find(filter: 'core.coderoot_set')! {
	// 	mut p := action.params
	// 	if p.exists('coderoot') {
	// 		coderoot := p.get_path_create('coderoot')!
	// 		mut gs := session.context.gitstructure()!
	// 		if gs.rootpath.path != coderoot {
	// 			mut db := session.context.contextdb.db_get(dbname: 'context')!
	// 			db.set('coderoot', coderoot)!
	// 			session.context.gitstructure_reload()!
	// 		}
	// 	} else {
	// 		return error('coderoot needs to be specified')
	// 	}
	// 	action.done = true
	// }

	// for mut action in plbook.find(filter: 'core.params_context_set')! {
	// 	mut p := action.params
	// 	for param in p.params {
	// 		session.context.params.set(param.key, param.value)
	// 	}
	// 	action.done = true
	// }

	// for mut action in plbook.find(filter: 'core.params_session_set')! {
	// 	mut p := action.params
	// 	for param in p.params {
	// 		session.params.set(param.key, param.value)
	// 	}
	// 	action.done = true
	// }

}
