module mcp
