module main

import freeflowuniverse.herolib.threefold.deploy

fn main() {
}
