module generic

// import freeflowuniverse.herolib.ui.console
// import freeflowuniverse.herolib.ui.telegram { UITelegram }
import freeflowuniverse.herolib.ui.uimodel

// ...
// ```
// args:
// TODO
// }
// ```
pub fn (mut c UserInterface) pay(args uimodel.PayArgs) ! {
	// match mut c.channel {
	// 	UIConsole { return c.channel.editor(args)! }
	// 	else { panic("can't find channel") }
	// }
}
