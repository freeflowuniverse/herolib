module code


pub type Value = string
