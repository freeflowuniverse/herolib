
module zerodb_client

import freeflowuniverse.herolib.core.base
import freeflowuniverse.herolib.core.playbook
import freeflowuniverse.herolib.ui.console


__global (
    zerodb_client_global map[string]&ZeroDBClient
    zerodb_client_default string
)

/////////FACTORY






