module currency

pub fn refresh() ! {
	d := {
		'USDAED': 3.673042
		'USDAFN': 67.503991
		'USDALL': 90.350403
		'USDAMD': 387.170403
		'USDANG': 1.803359
		'USDAOA': 912.503981
		'USDARS': 973.490388
		'USDAUD': 1.481262
		'USDAWG': 1.8005
		'USDAZN': 1.70397
		'USDBAM': 1.789575
		'USDBBD': 2.020322
		'USDBDT': 119.573423
		'USDBGN': 1.78838
		'USDBHD': 0.376903
		'USDBIF': 2893.5
		'USDBMD': 1
		'USDBND': 1.306987
		'USDBOB': 6.939367
		'USDBRL': 5.611304
		'USDBSD': 1.000645
		'USDBTC': 1.5975459e-5
		'USDBTN': 84.092851
		'USDBWP': 13.279045
		'USDBYN': 3.274501
		'USDBYR': 19600
		'USDBZD': 2.016881
		'USDCAD': 1.37705
		'USDCDF': 2878.000362
		'USDCHF': 0.857219
		'USDCLF': 0.033584
		'USDCLP': 926.680396
		'USDCNY': 7.066204
		'USDCNH': 7.073041
		'USDCOP': 4210.29
		'USDCRC': 516.884056
		'USDCUC': 1
		'USDCUP': 26.5
		'USDCVE': 101.290394
		'USDCZK': 23.126804
		'USDDJF': 177.720393
		'USDDKK': 6.821304
		'USDDOP': 60.40504
		'USDDZD': 132.93575
		'USDEGP': 48.517284
		'USDERN': 15
		'USDETB': 121.39275
		'USDEUR': 0.91335
		'USDFJD': 2.230391
		'USDFKP': 0.761559
		'USDGBP': 0.765169
		'USDGEL': 2.71504
		'USDGGP': 0.761559
		'USDGHS': 15.95504
		'USDGIP': 0.761559
		'USDGMD': 68.503851
		'USDGNF': 8636.000355
		'USDGTQ': 7.736965
		'USDGYD': 209.343075
		'USDHKD': 7.76988
		'USDHNL': 24.91504
		'USDHRK': 6.799011
		'USDHTG': 131.833342
		'USDHUF': 366.890388
		'USDIDR': 15569.15
		'USDILS': 3.75883
		'USDIMP': 0.761559
		'USDINR': 84.13735
		'USDIQD': 1309.5
		'USDIRR': 42102.503816
		'USDISK': 136.650386
		'USDJEP': 0.761559
		'USDJMD': 158.41557
		'USDJOD': 0.708504
		'USDJPY': 149.13904
		'USDKES': 129.000351
		'USDKGS': 85.503799
		'USDKHR': 4065.00035
		'USDKMF': 449.503794
		'USDKPW': 899.999433
		'USDKRW': 1349.320383
		'USDKWD': 0.30653
		'USDKYD': 0.833818
		'USDKZT': 484.459206
		'USDLAK': 21880.000349
		'USDLBP': 89600.000349
		'USDLKR': 292.894495
		'USDLRD': 192.803772
		'USDLSL': 17.490381
		'USDLTL': 2.95274
		'USDLVL': 0.60489
		'USDLYD': 4.795039
		'USDMAD': 9.803504
		'USDMDL': 17.659949
		'USDMGA': 4585.000347
		'USDMKD': 56.373726
		'USDMMK': 3247.960992
		'USDMNT': 3397.999955
		'USDMOP': 8.008821
		'USDMRU': 39.750379
		'USDMUR': 46.103741
		'USDMVR': 15.350378
		'USDMWK': 1736.000345
		'USDMXN': 19.279335
		'USDMYR': 4.287504
		'USDMZN': 63.903729
		'USDNAD': 17.490377
		'USDNGN': 1640.000344
		'USDNIO': 36.803722
		'USDNOK': 10.696745
		'USDNPR': 134.551493
		'USDNZD': 1.636822
		'USDOMR': 0.384447
		'USDPAB': 1.000618
		'USDPEN': 3.754604
		'USDPGK': 3.93225
		'USDPHP': 57.230375
		'USDPKR': 277.750374
		'USDPLN': 3.922272
		'USDPYG': 7809.426211
		'USDQAR': 3.641104
		'USDRON': 4.548504
		'USDRSD': 106.892552
		'USDRUB': 95.676332
		'USDRWF': 1355
		'USDSAR': 3.755532
		'USDSBD': 8.299327
		'USDSCR': 13.582042
		'USDSDG': 601.503676
		'USDSEK': 10.371445
		'USDSGD': 1.305104
		'USDSHP': 0.761559
		'USDSLE': 22.847303
		'USDSLL': 20969.494858
		'USDSOS': 571.000338
		'USDSRD': 31.946504
		'USDSTD': 20697.981008
		'USDSVC': 8.755725
		'USDSYP': 2512.529936
		'USDSZL': 17.403651
		'USDTHB': 33.155038
		'USDTJS': 10.666441
		'USDTMT': 3.51
		'USDTND': 3.071038
		'USDTOP': 2.342104
		'USDTRY': 34.281704
		'USDTTD': 6.791866
		'USDTWD': 32.178804
		'USDTZS': 2725.000335
		'USDUAH': 41.204244
		'USDUGX': 3677.388953
		'USDUYU': 41.843378
		'USDUZS': 12800.000334
		'USDVEF': 3622552.534434
		'USDVES': 38.83528
		'USDVND': 24820
		'USDVUV': 118.722009
		'USDWST': 2.797463
		'USDXAF': 600.184825
		'USDXAG': 0.031696
		'USDXAU': 0.000376
		'USDXCD': 2.70255
		'USDXDR': 0.744353
		'USDXOF': 598.503595
		'USDXPF': 109.550363
		'USDYER': 250.350363
		'USDZAR': 17.409585
		'USDZMK': 9001.203587
		'USDZMW': 26.440783
		'USDZWL': 321.999592
	}
	mut result := map[string]f64{}
	for name, val in d {
		name2 := name.all_after('USD')
		result[name2] = val
	}

	result['TFT'] = 0.01
	result['XLM'] = 0.092
	result['USDC'] = 1
	result['USD'] = 1

	lock currencies {
		for name, val in result {
			currencies[name] = Currency{
				name:   name
				usdval: val
			}
		}
	}
}
