module qdrant
