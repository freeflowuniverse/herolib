module heroprompt

import freeflowuniverse.herolib.core.base
import freeflowuniverse.herolib.core.playbook { PlayBook }
import freeflowuniverse.herolib.ui.console
import json
import os
import time

__global (
	heroprompt_global  map[string]&Workspace
	heroprompt_default string
)

/////////FACTORY

@[params]
pub struct ArgsGet {
pub mut:
	name   string = 'default'
	path   string
	fromdb bool // will load from filesystem
	create bool // default will not create if not exist
}

pub fn new(args ArgsGet) !&Workspace {
	// validate
	if args.name.len == 0 {
		return error('workspace name is required')
	}
	mut base_path := ''
	if args.path.len > 0 {
		if !os.exists(args.path) {
			return error('workspace path does not exist: ${args.path}')
		}
		if !os.is_dir(args.path) {
			return error('workspace path is not a directory: ${args.path}')
		}
		base_path = os.real_path(args.path)
	}
	mut obj := Workspace{
		name:      args.name
		base_path: base_path
		created:   time.now()
		updated:   time.now()
		is_saved:  false
	}
	set(obj)!
	return get(name: args.name)!
}

pub fn get(args ArgsGet) !&Workspace {
	mut context := base.context()!
	heroprompt_default = args.name
	if args.fromdb || args.name !in heroprompt_global {
		mut r := context.redis()!
		if r.hexists('context:heroprompt', args.name)! {
			data := r.hget('context:heroprompt', args.name)!
			if data.len == 0 {
				return error('Workspace with name: ${args.name} does not exist, prob bug.')
			}
			mut obj := json.decode(Workspace, data)!
			set_in_mem(obj)!
		} else {
			if args.create {
				new(args)!
			} else {
				return error("Workspace with name '${args.name}' does not exist")
			}
		}
		return get(name: args.name)! // no longer from db nor create
	}
	return heroprompt_global[args.name] or {
		return error('could not get config for heroprompt with name:heroprompt')
	}
}

// register the config for the future
pub fn set(o Workspace) ! {
	mut o2 := set_in_mem(o)!
	heroprompt_default = o2.name
	mut context := base.context()!
	mut r := context.redis()!
	r.hset('context:heroprompt', o2.name, json.encode(o2))!
}

// does the config exists?
pub fn exists(args ArgsGet) !bool {
	mut context := base.context()!
	mut r := context.redis()!
	return r.hexists('context:heroprompt', args.name)!
}

pub fn delete(args ArgsGet) ! {
	mut context := base.context()!
	mut r := context.redis()!
	r.hdel('context:heroprompt', args.name)!
}

@[params]
pub struct ArgsList {
pub mut:
	fromdb bool // will load from filesystem
}

// if fromdb set: load from filesystem, and not from mem, will also reset what is in mem
pub fn list(args ArgsList) ![]&Workspace {
	mut res := []&Workspace{}
	mut context := base.context()!
	if args.fromdb {
		// reset what is in mem
		heroprompt_global = map[string]&Workspace{}
		heroprompt_default = ''
	}
	if args.fromdb {
		mut r := context.redis()!
		mut l := r.hkeys('context:heroprompt')!

		for name in l {
			res << get(name: name, fromdb: true)!
		}
		return res
	} else {
		// load from memory
		for _, client in heroprompt_global {
			res << client
		}
	}
	return res
}

// only sets in mem, does not set as config
fn set_in_mem(o Workspace) !Workspace {
	mut o2 := obj_init(o)!
	heroprompt_global[o2.name] = &o2
	heroprompt_default = o2.name
	return o2
}

pub fn play(mut plbook PlayBook) ! {
	if !plbook.exists(filter: 'heroprompt.') {
		return
	}
	mut install_actions := plbook.find(filter: 'heroprompt.configure')!
	if install_actions.len > 0 {
		for install_action in install_actions {
			heroscript := install_action.heroscript()
			mut obj2 := heroscript_loads(heroscript)!
			set(obj2)!
		}
	}
}

// switch instance to be used for heroprompt
pub fn switch(name string) {
	heroprompt_default = name
}
