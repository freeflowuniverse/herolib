module datamodel

pub struct NodeSim {
	Node
pub mut:
	cost f64 // free
}
