module wireguard

fn (wg WireGuard) show() {
}

fn (wg WireGuard) up() {
}

fn (wg WireGuard) down() {
}

fn (wg WireGuard) generate_key() !string {
}

fn (wg WireGuard) get_public_key() {
}
