module rhai
