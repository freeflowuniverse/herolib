module datamodel
import freeflowuniverse.herolib.threefold.grid4.datamodel { Node }
pub struct NodeSim {
	Node
pub mut:
	cost f64 // free
}
