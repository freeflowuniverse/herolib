module models

import freeflowuniverse.herolib.data.encoder

// Standalone tests for the Wallet model that don't depend on other models

fn test_wallet_standalone_dumps_loads() {
	// Create a test wallet with sample data
	mut wallet := Wallet{
		id: 123
		name: 'Test Wallet'
		description: 'A test wallet for binary encoding'
		blockchain_name: 'Ethereum'
		pubkey: '0x123456789abcdef'
	}
	
	// Add assets
	wallet.assets << Asset{
		name: 'ETH'
		amount: 1.5
	}
	
	wallet.assets << Asset{
		name: 'USDC'
		amount: 1000.0
	}
	
	// Test binary encoding
	binary_data := wallet.dumps() or {
		assert false, 'Failed to encode wallet: ${err}'
		return
	}
	
	// Test binary decoding
	decoded_wallet := wallet_loads(binary_data) or {
		assert false, 'Failed to decode wallet: ${err}'
		return
	}
	
	// Verify the decoded data matches the original
	assert decoded_wallet.id == wallet.id
	assert decoded_wallet.name == wallet.name
	assert decoded_wallet.description == wallet.description
	assert decoded_wallet.blockchain_name == wallet.blockchain_name
	assert decoded_wallet.pubkey == wallet.pubkey
	
	// Verify assets
	assert decoded_wallet.assets.len == wallet.assets.len
	
	// Verify first asset
	assert decoded_wallet.assets[0].name == wallet.assets[0].name
	assert decoded_wallet.assets[0].amount == wallet.assets[0].amount
	
	// Verify second asset
	assert decoded_wallet.assets[1].name == wallet.assets[1].name
	assert decoded_wallet.assets[1].amount == wallet.assets[1].amount
	
	println('Wallet binary encoding/decoding test passed successfully')
}

fn test_wallet_standalone_set_asset() {
	mut wallet := Wallet{
		id: 456
		name: 'Asset Test Wallet'
		blockchain_name: 'Bitcoin'
		pubkey: 'bc1q123456789'
	}
	
	// Test adding a new asset
	wallet.set_asset('BTC', 0.5)
	assert wallet.assets.len == 1
	assert wallet.assets[0].name == 'BTC'
	assert wallet.assets[0].amount == 0.5
	
	// Test updating an existing asset
	wallet.set_asset('BTC', 1.0)
	assert wallet.assets.len == 1 // Should still have only one asset
	assert wallet.assets[0].name == 'BTC'
	assert wallet.assets[0].amount == 1.0 // Amount should be updated
	
	// Add another asset
	wallet.set_asset('USDT', 500.0)
	assert wallet.assets.len == 2
	
	// Verify both assets are present with correct values
	for asset in wallet.assets {
		if asset.name == 'BTC' {
			assert asset.amount == 1.0
		} else if asset.name == 'USDT' {
			assert asset.amount == 500.0
		} else {
			assert false, 'Unexpected asset: ${asset.name}'
		}
	}
	
	println('Wallet set_asset test passed successfully')
}

fn test_wallet_standalone_total_value() {
	mut wallet := Wallet{
		id: 789
		name: 'Value Test Wallet'
		blockchain_name: 'Solana'
		pubkey: 'sol123456789'
	}
	
	// Empty wallet should have zero value
	assert wallet.total_value() == 0.0
	
	// Add first asset
	wallet.set_asset('SOL', 10.0)
	assert wallet.total_value() == 10.0
	
	// Add second asset
	wallet.set_asset('USDC', 50.0)
	assert wallet.total_value() == 60.0 // 10 SOL + 50 USDC
	
	// Update first asset
	wallet.set_asset('SOL', 15.0)
	assert wallet.total_value() == 65.0 // 15 SOL + 50 USDC
	
	// Add third asset with negative value
	wallet.set_asset('TEST', -5.0)
	assert wallet.total_value() == 60.0 // 15 SOL + 50 USDC - 5 TEST
	
	println('Wallet total_value test passed successfully')
}

fn test_wallet_standalone_index_keys() {
	wallet := Wallet{
		id: 101
		name: 'Index Keys Test'
		blockchain_name: 'Polkadot'
		pubkey: 'dot123456789'
	}
	
	keys := wallet.index_keys()
	assert keys['name'] == 'Index Keys Test'
	assert keys['blockchain'] == 'Polkadot'
	assert keys.len == 2
	
	println('Wallet index_keys test passed successfully')
}

fn test_wallet_standalone_wrong_encoding_id() {
	// Create invalid data with wrong encoding ID
	mut e := encoder.new()
	e.add_u16(999) // Wrong ID (should be 202)
	
	// Attempt to deserialize and expect error
	result := wallet_loads(e.data) or {
		assert err.str() == 'Wrong file type: expected encoding ID 202, got 999, for wallet'
		println('Error handling test (wrong encoding ID) passed successfully')
		return
	}
	
	assert false, 'Should have returned an error for wrong encoding ID'
}

fn main() {
	test_wallet_standalone_dumps_loads()
	test_wallet_standalone_set_asset()
	test_wallet_standalone_total_value()
	test_wallet_standalone_index_keys()
	test_wallet_standalone_wrong_encoding_id()
	
	println('All Wallet standalone tests passed successfully')
}