module gitea_client
