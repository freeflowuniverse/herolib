module stage

