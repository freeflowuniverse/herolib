module docusaurus

import freeflowuniverse.herolib.develop.gittools
import freeflowuniverse.herolib.osal
import freeflowuniverse.herolib.installers.web.bun
import freeflowuniverse.herolib.core.pathlib
import json
import os
import time

@[params]
struct TemplateInstallArgs {
	template_update bool = true
	install         bool
	delete          bool = true
}

fn (mut self DocusaurusFactory) template_install(args TemplateInstallArgs) ! {
	mut gs := gittools.new()!

	mut r := gs.get_repo(
		url:  'https://github.com/freeflowuniverse/docusaurus_template.git'
		pull: args.template_update
	)!
	mut template_path := r.patho()!

	// always start from template first for static assets and source files
	for item in ['src', 'static'] {
		mut aa := template_path.dir_get(item)!
		aa.copy(dest: '${self.path_build.path}/${item}', delete: args.delete)!
	}

	// Generate config files dynamically from config
	self.generate_package_json()!
	self.generate_tsconfig_json()!
	self.generate_sidebars_ts()!
	self.generate_docusaurus_config_ts()!

	if args.install {
		// install bun
		mut installer := bun.get()!
		installer.install()!

		osal.exec(
			cmd: '
				${osal.profile_path_source_and()!} 
				export PATH=/tmp/docusaurus_build/node_modules/.bin:${os.home_dir()}/.bun/bin/:??PATH
				cd ${self.path_build.path}
				bun install
			'
		)!
	}

	// Only try to delete docs if it exists in the template
	if os.exists(os.join_path(template_path.path, 'docs')) {
		mut aa := template_path.dir_get('docs')!
		aa.delete()!
	}
}

// Generate package.json based on the configuration
fn (mut self DocusaurusFactory) generate_package_json() ! {
	// Build package.json content as a structured JSON string
	mut name := 'docusaurus-site'
	if self.config.main.name != '' {
		name = self.config.main.name
	} else if self.config.navbar.title != '' {
		name = self.config.navbar.title.to_lower().replace(' ', '-')
	}

	// Create the JSON structure manually
	package_json := '{
	 "name": "${name}",
	 "version": "0.0.1",
	 "private": true,
	 "scripts": {
	   "docusaurus": "docusaurus",
	   "start": "docusaurus start",
	   "build": "docusaurus build",
	   "swizzle": "docusaurus swizzle",
	   "deploy": "docusaurus deploy",
	   "clear": "docusaurus clear",
	   "serve": "docusaurus serve",
	   "write-translations": "docusaurus write-translations",
	   "write-heading-ids": "docusaurus write-heading-ids",
	   "typecheck": "tsc"
	 },
	 "dependencies": {
	   "@docusaurus/core": "^3.1.0",
	   "@docusaurus/preset-classic": "^3.1.0",
	   "@mdx-js/react": "^3.0.0",
	   "clsx": "^2.0.0",
	   "prism-react-renderer": "^2.3.0",
	   "react": "^18.0.0",
	   "react-dom": "^18.0.0"
	 },
	 "devDependencies": {
	   "@docusaurus/module-type-aliases": "^3.1.0",
	   "@docusaurus/tsconfig": "^3.1.0",
	   "@docusaurus/types": "^3.1.0",
	   "typescript": "^5.2.2"
	 },
	 "browserslist": {
	   "production": [">0.5%", "not dead", "not op_mini all"],
	   "development": ["last 1 chrome version", "last 1 firefox version", "last 1 safari version"]
	 },
	 "engines": {
	   "node": ">=18.0"
	 }
}' // Write to file

	mut package_file := pathlib.get_file(
		path:   os.join_path(self.path_build.path, 'package.json')
		create: true
	)!
	package_file.write(package_json)!
}

// Generate tsconfig.json based on the configuration
fn (mut self DocusaurusFactory) generate_tsconfig_json() ! {
	// Create tsconfig.json as a manual JSON string
	tsconfig_json := '{
	 "extends": "@docusaurus/tsconfig",
	 "compilerOptions": {
	   "baseUrl": ".",
	   "resolveJsonModule": true
	 },
	 "include": ["src/**/*", "docusaurus.config.ts"]
}'

	// Write to file
	mut tsconfig_file := pathlib.get_file(
		path:   os.join_path(self.path_build.path, 'tsconfig.json')
		create: true
	)!
	tsconfig_file.write(tsconfig_json)!
}

// Generate sidebars.ts based on the configuration
fn (mut self DocusaurusFactory) generate_sidebars_ts() ! {
	// Simple default sidebar structure
	sidebar_content := "import type {SidebarsConfig} from '@docusaurus/plugin-content-docs';

/**
	* Creating a sidebar enables you to:
	- create an ordered group of docs
	- render a sidebar for each doc of that group
	- provide next/previous navigation

	The sidebars can be generated from the filesystem, or explicitly defined here.

	Create as many sidebars as you want.
	*/
const sidebars: SidebarsConfig = {
	 // By default, Docusaurus generates a sidebar from the docs folder structure
	 tutorialSidebar: [{type: 'autogenerated', dirName: '.'}],
};

export default sidebars;
"
	mut sidebars_file := pathlib.get_file(
		path:   os.join_path(self.path_build.path, 'sidebars.ts')
		create: true
	)!
	sidebars_file.write(sidebar_content)!
}

// Generate docusaurus.config.ts based on the configuration
fn (mut self DocusaurusFactory) generate_docusaurus_config_ts() ! {
	// Use config values with fallbacks
	title := if self.config.main.title != '' { self.config.main.title } else { 'Docusaurus Site' }
	tagline := if self.config.main.tagline != '' {
		self.config.main.tagline
	} else {
		'Documentation Site'
	}
	url := if self.config.main.url != '' { self.config.main.url } else { 'https://example.com' }
	base_url := if self.config.main.base_url != '' { self.config.main.base_url } else { '/' }
	favicon := if self.config.main.favicon != '' {
		self.config.main.favicon
	} else {
		'img/favicon.png'
	}

	// Format navbar items from config
	mut navbar_items := []string{}
	for item in self.config.navbar.items {
		navbar_items << "{
			label: '${item.label}',
			href: '${item.href}',
			position: '${item.position}'
		}"
	}

	navbar_items_str := navbar_items.join(',\n      ')

	// Generate footer links if available
	mut footer_links := []string{}
	for link in self.config.footer.links {
		mut items := []string{}
		for item in link.items {
			mut item_str := '{'
			if item.label != '' {
				item_str += "label: '${item.label}', "
			}

			// Ensure only one of 'to', 'href', or 'html' is used
			// Priority: href > to > html
			if item.href != '' {
				item_str += "href: '${item.href}'"
			} else if item.to != '' {
				item_str += "to: '${item.to}'"
			} else {
				// Default to linking to docs if nothing specified
				item_str += "to: '/docs'"
			}

			item_str += '}'
			items << item_str
		}

		footer_links << "{
			title: '${link.title}',
			items: [
				${items.join(',\n          ')}
			]
		}"
	}

	footer_links_str := footer_links.join(',\n      ')

	// Year for copyright
	year := time.now().year.str()

	copyright := if self.config.main.copyright != '' {
		self.config.main.copyright
	} else {
		'Copyright © ${year} ${title}'
	}

	// Construct the full config file content
	config_content := "import {themes as prismThemes} from 'prism-react-renderer';
import type {Config} from '@docusaurus/types';
import type * as Preset from '@docusaurus/preset-classic';

const config: Config = {
	 title: '${title}',
	 tagline: '${tagline}',
	 favicon: '${favicon}',
	 
	 // Set the production url of your site here
	 url: '${url}',
	 // Set the /<baseUrl>/ pathname under which your site is served
	 // For GitHub pages deployment, it is often '/<projectName>/'
	 baseUrl: '${base_url}',

	 // GitHub pages deployment config.
	 // If you aren't using GitHub pages, you don't need these.
	 organizationName: 'freeflowuniverse', // Usually your GitHub org/user name.
	 projectName: '${self.config.main.name}', // Usually your repo name.

	 onBrokenLinks: 'warn',
	 onBrokenMarkdownLinks: 'warn',
	 
	 // Enable for i18n
	 // i18n: {
	 //   defaultLocale: 'en',
	 //   locales: ['en'],
	 // },

	 presets: [
	   [
	     'classic',
	     {
	       docs: {
	         sidebarPath: './sidebars.ts',
	       },
	       theme: {
	         customCss: './src/css/custom.css',
	       },
	     } satisfies Preset.Options,
	   ],
	 ],

	 themeConfig: {
	   // Replace with your project's social card
	   image: 'img/docusaurus-social-card.jpg',
	   navbar: {
	     title: '${self.config.navbar.title}',
	     logo: {
	       alt: 'Logo',
	       src: 'img/logo.svg',
	     },
	     items: [
	       ${navbar_items_str}
	     ],
	   },
	   footer: {
	     style: '${self.config.footer.style}',
	     links: [
	       ${footer_links_str}
	     ],
	     copyright: '${copyright}',
	   },
	   prism: {
	     theme: prismThemes.github,
	     darkTheme: prismThemes.dracula,
	   },
	 } satisfies Preset.ThemeConfig,
};

export default config;
"

	mut config_file := pathlib.get_file(
		path:   os.join_path(self.path_build.path, 'docusaurus.config.ts')
		create: true
	)!
	config_file.write(config_content)!
}
