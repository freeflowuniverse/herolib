module cloudslices




