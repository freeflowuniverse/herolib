module ourdb

fn test_basic_operations() {
	// mut client := get()
}
