module streamer
