module gitea_client

//PUT the models for swagger here