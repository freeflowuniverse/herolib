module template

// import os
import freeflowuniverse.herolib.ui.uimodel { QuestionArgs }
// import freeflowuniverse.herolib.ui.console

// args:
// - description string
// - question string
// - warning: string (if it goes wrong, which message to use)
// - reset bool = true
// - regex: to check what result need to be part of
// - minlen: min nr of chars
//
pub fn (mut c UIExample) ask_question(args QuestionArgs) !string {
	return ''
}
