module python

import freeflowuniverse.herolib.data.encoderhero

pub const version = '3.12.0'
const singleton = true
const default = true

// THIS THE THE SOURCE OF THE INFORMATION OF THIS FILE, HERE WE HAVE THE CONFIG OBJECT CONFIGURED AND MODELLED
@[heap]
pub struct Python {
pub mut:
	name string = 'default'
}

// your checking & initialization code if needed
fn obj_init(mycfg_ Python) !Python {
	mut mycfg := mycfg_
	return mycfg
}

// called before start if done
fn configure() ! {
	// mut installer := get()!
}

/////////////NORMALLY NO NEED TO TOUCH

pub fn heroscript_dumps(obj Python) !string {
	return encoderhero.encode[Python](obj)!
}

pub fn heroscript_loads(heroscript string) !Python {
	mut obj := encoderhero.decode[Python](heroscript)!
	return obj
}
