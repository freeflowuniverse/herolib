module developer

pub struct Developer {}

