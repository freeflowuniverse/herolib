module developer

import freeflowuniverse.herolib.mcp

// Tool definition for the create_mcp_tool function
const create_mcp_tool_tool = mcp.Tool{
	name: 'create_mcp_tool'
	description: 'Parses a V language function string and returns an MCP Tool struct. This tool analyzes function signatures, extracts parameters, and generates the appropriate MCP Tool representation.'
	input_schema: mcp.ToolInputSchema{
		typ: 'object'
		properties: {
			'function': mcp.ToolProperty{
				typ: 'string'
			}
			'types': mcp.ToolProperty{
				typ: 'object'
			}
		}
		required: ['function']
	}
}
