module codewalker

pub struct Error {
pub:
	message string
	linenr  int
	category string
}