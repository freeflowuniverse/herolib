module stage
