module mycelium

